----------------------------------------------------------------------
-- ¡IMPORTANTE! Rellene la cabecera del fichero
-- Fecha:
-- Autores:
----------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

entity ExtCero is
    port ( 
		A : IN  unsigned(7 downto 0);
		Q : OUT  unsigned(11 downto 0)
	);
end ExtCero;

architecture Practica of ExtCero is

begin
	
end Practica;
